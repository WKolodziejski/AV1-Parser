library ieee;
use ieee.std_logic_1164.all;
        use IEEE.std_logic_signed.all;

use ieee.numeric_std.all; 
--use ieee.std_logic_arith.all;


entity Escolha is
	port(vet_sel: in std_logic_vector(7 downto 0);
		  S0, S3: out std_logic_vector(2 downto 0);
		  S1, S2: out std_logic_vector(5 downto 0);
		  sinalA0, sinalA1: out std_logic
        );
end Escolha;


architecture comportamento of Escolha is
	signal aux8: signed (1 downto 0);
	begin 
	process (vet_sel)
	begin

		case vet_sel is

------------------------- Filtro 1------------------------------

			when "00000000" => --[0, 128, 0, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "001001";
				S2 <= "001001";
				S3 <= "000";
				sinalA1 <= '0';

			when "00000001" => --[8, 108, 8, 4]
				S0 <= "011";
				sinalA0 <= '0';
				S1 <= "000111";
				S2 <= "000000";
				S3 <= "010";
				sinalA1 <= '0';

			when "00000010" => --[-4, 108, 16, 8]
				S0 <= "010";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000001";
				S3 <= "011";
				sinalA1 <= '1';

			when "00000011" => --[-8, 108, 32, -4]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000011";
				S3 <= "010";
				sinalA1 <= '1';

			when "00000100" => --[-8, 108, 44, -16]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000100";
				S3 <= "100";
				sinalA1 <= '1';

			when "00000101" => --[-16, 108, 44, -8]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000100";
				S3 <= "011";
				sinalA1 <= '1';

			when "00000110" => --[-16, 84, 64, -4]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000110";
				S2 <= "000101";
				S3 <= "010";
				sinalA1 <= '1';

			when "00000111" => --[-16, 84, 64, -4]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000110";
				S2 <= "000101";
				S3 <= "010";
				sinalA1 <= '1';

			when "00001000" => --[-32, 84, 84, -8]
				S0 <= "101";
				sinalA0 <= '1';
				S1 <= "000110";
				S2 <= "000110";
				S3 <= "011";
				sinalA1 <= '1';

			when "00001001" => --[-4, 64, 84, -16]
				S0 <= "010";
				sinalA0 <= '1';
				S1 <= "000101";
				S2 <= "000110";
				S3 <= "100";
				sinalA1 <= '1';

			when "00001010" => --[-4, 64, 84, -16]
				S0 <= "010";
				sinalA0 <= '1';
				S1 <= "000101";
				S2 <= "000110";
				S3 <= "100";
				sinalA1 <= '1';

			when "00001011" => --[-8, 44, 108, -16]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000100";
				S2 <= "000111";
				S3 <= "100";
				sinalA1 <= '1';

			when "00001100" => --[-16, 44, 108, -8]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000100";
				S2 <= "000111";
				S3 <= "011";
				sinalA1 <= '1';

			when "00001101" => --[-4, 32, 108, -8]
				S0 <= "010";
				sinalA0 <= '1';
				S1 <= "000011";
				S2 <= "000111";
				S3 <= "011";
				sinalA1 <= '1';

			when "00001110" => --[8, 16, 108, -4]
				S0 <= "011";
				sinalA0 <= '0';
				S1 <= "000001";
				S2 <= "000111";
				S3 <= "010";
				sinalA1 <= '0';

			when "00001111" => --[4, 8, 108, 8]
				S0 <= "010";
				sinalA0 <= '0';
				S1 <= "000000";
				S2 <= "000111";
				S3 <= "011";
				sinalA1 <= '0';

------------------------- Filtro 2------------------------------

			when "00010000" => --[0, 128, 0, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "001001";
				S2 <= "001001";
				S3 <= "000";
				sinalA1 <= '0';

			when "00010001" => --[32, 64, 32, 0]
				S0 <= "101";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000011";
				S3 <= "000";
				sinalA1 <= '0';

			when "00010010" => --[32, 64, 32, 0]
				S0 <= "101";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000011";
				S3 <= "000";
				sinalA1 <= '0';

			when "00010011" => --[32, 64, 32, 0]
				S0 <= "101";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000011";
				S3 <= "000";
				sinalA1 <= '0';

			when "00010100" => --[32, 64, 32, 0]
				S0 <= "101";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000011";
				S3 <= "000";
				sinalA1 <= '0';

			when "00010101" => --[16, 64, 32, 16]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000011";
				S3 <= "100";
				sinalA1 <= '0';

			when "00010110" => --[16, 64, 32, 16]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000011";
				S3 <= "100";
				sinalA1 <= '0';

			when "00010111" => --[16, 64, 32, 16]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000011";
				S3 <= "100";
				sinalA1 <= '0';

			when "00011000" => --[32, 44, 44, 8]
				S0 <= "101";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000100";
				S3 <= "011";
				sinalA1 <= '0';

			when "00011001" => --[16, 32, 64, 16]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000011";
				S2 <= "000101";
				S3 <= "100";
				sinalA1 <= '0';

			when "00011010" => --[16, 32, 64, 16]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000011";
				S2 <= "000101";
				S3 <= "100";
				sinalA1 <= '0';

			when "00011011" => --[16, 32, 64, 16]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000011";
				S2 <= "000101";
				S3 <= "100";
				sinalA1 <= '0';

			when "00011100" => --[0, 32, 64, 32]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000011";
				S2 <= "000101";
				S3 <= "101";
				sinalA1 <= '0';

			when "00011101" => --[0, 32, 64, 32]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000011";
				S2 <= "000101";
				S3 <= "101";
				sinalA1 <= '0';

			when "00011110" => --[0, 32, 64, 32]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000011";
				S2 <= "000101";
				S3 <= "101";
				sinalA1 <= '0';

			when "00011111" => --[0, 32, 64, 32]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000011";
				S2 <= "000101";
				S3 <= "101";
				sinalA1 <= '0';

------------------------- Filtro 3------------------------------

			when "00100000" => --[0, 128, 0, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "001001";
				S2 <= "001001";
				S3 <= "000";
				sinalA1 <= '0';

			when "00100001" => --[4, 108, 8, 8]
				S0 <= "010";
				sinalA0 <= '0';
				S1 <= "000111";
				S2 <= "000000";
				S3 <= "011";
				sinalA1 <= '0';

			when "00100010" => --[-8, 108, 32, -4]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000011";
				S3 <= "010";
				sinalA1 <= '1';

			when "00100011" => --[-8, 108, 32, -4]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000011";
				S3 <= "010";
				sinalA1 <= '1';

			when "00100100" => --[-16, 108, 44, -8]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000100";
				S3 <= "011";
				sinalA1 <= '1';

			when "00100101" => --[-16, 108, 44, -8]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000100";
				S3 <= "011";
				sinalA1 <= '1';

			when "00100110" => --[-32, 108, 64, -16]
				S0 <= "101";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000101";
				S3 <= "100";
				sinalA1 <= '1';

			when "00100111" => --[-32, 84, 84, -8]
				S0 <= "101";
				sinalA0 <= '1';
				S1 <= "000110";
				S2 <= "000110";
				S3 <= "011";
				sinalA1 <= '1';

			when "00101000" => --[-32, 84, 84, -8]
				S0 <= "101";
				sinalA0 <= '1';
				S1 <= "000110";
				S2 <= "000110";
				S3 <= "011";
				sinalA1 <= '1';

			when "00101001" => --[-8, 84, 84, -32]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000110";
				S2 <= "000110";
				S3 <= "101";
				sinalA1 <= '1';

			when "00101010" => --[-16, 64, 108, -32]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000101";
				S2 <= "000111";
				S3 <= "101";
				sinalA1 <= '1';

			when "00101011" => --[-8, 44, 108, -16]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000100";
				S2 <= "000111";
				S3 <= "100";
				sinalA1 <= '1';

			when "00101100" => --[-8, 44, 108, -16]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000100";
				S2 <= "000111";
				S3 <= "100";
				sinalA1 <= '1';

			when "00101101" => --[-4, 32, 108, -8]
				S0 <= "010";
				sinalA0 <= '1';
				S1 <= "000011";
				S2 <= "000111";
				S3 <= "011";
				sinalA1 <= '1';

			when "00101110" => --[-4, 32, 108, -8]
				S0 <= "010";
				sinalA0 <= '1';
				S1 <= "000011";
				S2 <= "000111";
				S3 <= "011";
				sinalA1 <= '1';

			when "00101111" => --[8, 8, 108, 4]
				S0 <= "011";
				sinalA0 <= '0';
				S1 <= "000000";
				S2 <= "000111";
				S3 <= "010";
				sinalA1 <= '0';

------------------------- Filtro 4------------------------------

			when "00110000" => --[0, 128, 0, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "001001";
				S2 <= "001001";
				S3 <= "000";
				sinalA1 <= '0';

			when "00110001" => --[0, 108, 20, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000111";
				S2 <= "000010";
				S3 <= "000";
				sinalA1 <= '0';

			when "00110010" => --[0, 108, 20, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000111";
				S2 <= "000010";
				S3 <= "000";
				sinalA1 <= '0';

			when "00110011" => --[0, 108, 20, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000111";
				S2 <= "000010";
				S3 <= "000";
				sinalA1 <= '0';

			when "00110100" => --[0, 108, 20, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000111";
				S2 <= "000010";
				S3 <= "000";
				sinalA1 <= '0';

			when "00110101" => --[0, 84, 44, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000110";
				S2 <= "000100";
				S3 <= "000";
				sinalA1 <= '0';

			when "00110110" => --[0, 84, 44, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000110";
				S2 <= "000100";
				S3 <= "000";
				sinalA1 <= '0';

			when "00110111" => --[0, 84, 44, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000110";
				S2 <= "000100";
				S3 <= "000";
				sinalA1 <= '0';

			when "00111000" => --[0, 64, 64, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000101";
				S3 <= "000";
				sinalA1 <= '0';

			when "00111001" => --[0, 44, 84, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000110";
				S3 <= "000";
				sinalA1 <= '0';

			when "00111010" => --[0, 44, 84, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000110";
				S3 <= "000";
				sinalA1 <= '0';

			when "00111011" => --[0, 44, 84, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000110";
				S3 <= "000";
				sinalA1 <= '0';

			when "00111100" => --[0, 20, 108, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000010";
				S2 <= "000111";
				S3 <= "000";
				sinalA1 <= '0';

			when "00111101" => --[0, 20, 108, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000010";
				S2 <= "000111";
				S3 <= "000";
				sinalA1 <= '0';

			when "00111110" => --[0, 20, 108, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000010";
				S2 <= "000111";
				S3 <= "000";
				sinalA1 <= '0';

			when "00111111" => --[0, 20, 108, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000010";
				S2 <= "000111";
				S3 <= "000";
				sinalA1 <= '0';

------------------------- Filtro 5------------------------------

			when "01000000" => --[0, 128, 0, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "001001";
				S2 <= "001001";
				S3 <= "000";
				sinalA1 <= '0';

			when "01000001" => --[8, 108, 8, 4]
				S0 <= "011";
				sinalA0 <= '0';
				S1 <= "000111";
				S2 <= "000000";
				S3 <= "010";
				sinalA1 <= '0';

			when "01000010" => --[2, 108, 16, 2]
				S0 <= "001";
				sinalA0 <= '0';
				S1 <= "000111";
				S2 <= "000001";
				S3 <= "001";
				sinalA1 <= '0';

			when "01000011" => --[-8, 108, 32, -4]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000011";
				S3 <= "010";
				sinalA1 <= '1';

			when "01000100" => --[-16, 108, 44, -8]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000100";
				S3 <= "011";
				sinalA1 <= '1';

			when "01000101" => --[-16, 108, 44, -8]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000111";
				S2 <= "000100";
				S3 <= "011";
				sinalA1 <= '1';

			when "01000110" => --[-16, 84, 64, -4]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000110";
				S2 <= "000101";
				S3 <= "010";
				sinalA1 <= '1';

			when "01000111" => --[-16, 84, 64, -4]
				S0 <= "100";
				sinalA0 <= '1';
				S1 <= "000110";
				S2 <= "000101";
				S3 <= "010";
				sinalA1 <= '1';

			when "01001000" => --[-32, 84, 84, -8]
				S0 <= "101";
				sinalA0 <= '1';
				S1 <= "000110";
				S2 <= "000110";
				S3 <= "011";
				sinalA1 <= '1';

			when "01001001" => --[-4, 64, 84, -16]
				S0 <= "010";
				sinalA0 <= '1';
				S1 <= "000101";
				S2 <= "000110";
				S3 <= "100";
				sinalA1 <= '1';

			when "01001010" => --[-4, 64, 84, -16]
				S0 <= "010";
				sinalA0 <= '1';
				S1 <= "000101";
				S2 <= "000110";
				S3 <= "100";
				sinalA1 <= '1';

			when "01001011" => --[-8, 44, 108, -16]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000100";
				S2 <= "000111";
				S3 <= "100";
				sinalA1 <= '1';

			when "01001100" => --[-8, 44, 108, -16]
				S0 <= "011";
				sinalA0 <= '1';
				S1 <= "000100";
				S2 <= "000111";
				S3 <= "100";
				sinalA1 <= '1';

			when "01001101" => --[-4, 32, 108, -8]
				S0 <= "010";
				sinalA0 <= '1';
				S1 <= "000011";
				S2 <= "000111";
				S3 <= "011";
				sinalA1 <= '1';

			when "01001110" => --[2, 16, 108, 2]
				S0 <= "001";
				sinalA0 <= '0';
				S1 <= "000001";
				S2 <= "000111";
				S3 <= "001";
				sinalA1 <= '0';

			when "01001111" => --[4, 8, 108, 8]
				S0 <= "010";
				sinalA0 <= '0';
				S1 <= "000000";
				S2 <= "000111";
				S3 <= "011";
				sinalA1 <= '0';

------------------------- Filtro 6------------------------------

			when "01010000" => --[0, 128, 0, 0]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "001001";
				S2 <= "001001";
				S3 <= "000";
				sinalA1 <= '0';

			when "01010001" => --[32, 64, 32, 0]
				S0 <= "101";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000011";
				S3 <= "000";
				sinalA1 <= '0';

			when "01010010" => --[32, 64, 32, 0]
				S0 <= "101";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000011";
				S3 <= "000";
				sinalA1 <= '0';

			when "01010011" => --[16, 64, 44, 4]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000100";
				S3 <= "010";
				sinalA1 <= '0';

			when "01010100" => --[16, 64, 44, 4]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000100";
				S3 <= "010";
				sinalA1 <= '0';

			when "01010101" => --[16, 64, 44, 4]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000100";
				S3 <= "010";
				sinalA1 <= '0';

			when "01010110" => --[16, 64, 44, 4]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000100";
				S3 <= "010";
				sinalA1 <= '0';

			when "01010111" => --[16, 64, 44, 4]
				S0 <= "100";
				sinalA0 <= '0';
				S1 <= "000101";
				S2 <= "000100";
				S3 <= "010";
				sinalA1 <= '0';

			when "01011000" => --[32, 44, 44, 8]
				S0 <= "101";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000100";
				S3 <= "011";
				sinalA1 <= '0';

			when "01011001" => --[4, 44, 64, 16]
				S0 <= "010";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000101";
				S3 <= "100";
				sinalA1 <= '0';

			when "01011010" => --[4, 44, 64, 16]
				S0 <= "010";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000101";
				S3 <= "100";
				sinalA1 <= '0';

			when "01011011" => --[4, 44, 64, 16]
				S0 <= "010";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000101";
				S3 <= "100";
				sinalA1 <= '0';

			when "01011100" => --[4, 44, 64, 16]
				S0 <= "010";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000101";
				S3 <= "100";
				sinalA1 <= '0';

			when "01011101" => --[4, 44, 64, 16]
				S0 <= "010";
				sinalA0 <= '0';
				S1 <= "000100";
				S2 <= "000101";
				S3 <= "100";
				sinalA1 <= '0';

			when "01011110" => --[0, 32, 64, 32]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000011";
				S2 <= "000101";
				S3 <= "101";
				sinalA1 <= '0';

			when "01011111" => --[0, 32, 64, 32]
				S0 <= "000";
				sinalA0 <= '0';
				S1 <= "000011";
				S2 <= "000101";
				S3 <= "101";
				sinalA1 <= '0';

			when others =>
				aux8 <= "00";
		
		end case;

	end process;

end comportamento;