library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_signed.all;
use ieee.numeric_std.all; 

entity Escolha is
	port(vet_sel: in std_logic_vector(7 downto 0);
		S0, S3: out std_logic_vector(2 downto 0);
		S1, S2: out std_logic_vector(5 downto 0);
		sinalA0, sinalA1: out std_logic
		);
end Escolha;


architecture comportamento of Escolha is
	signal aux8: signed (1 downto 0);
	begin
	process (vet_sel)
	begin

		case vet_sel is

------------------------- Filtro 1------------------------------

			when "00000000" => --[0, 0, 127, 1, 0, 0, 0, 0]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "01111111";
				S3 <= "00000001";
				S4 <= "00000000";
				S5 <= "00000000";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00000001" => --[0, -1, 127, 2, 0, 0, 0, 0]
				S0 <= "00000000";
				S1 <= "00000001";
				S2 <= "01111111";
				S3 <= "00000010";
				S4 <= "00000000";
				S5 <= "00000000";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00000010" => --[1, -3, 127, 4, -1, 0, 0, 0]
				S0 <= "00000001";
				S1 <= "00000011";
				S2 <= "01111111";
				S3 <= "00000100";
				S4 <= "00000001";
				S5 <= "00000000";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00000011" => --[1, -4, 126, 6, -2, 1, 0, 0]
				S0 <= "00000001";
				S1 <= "00000100";
				S2 <= "01111110";
				S3 <= "00000110";
				S4 <= "00000010";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00000100" => --[1, -5, 126, 8, -3, 1, 0, 0]
				S0 <= "00000001";
				S1 <= "00000101";
				S2 <= "01111110";
				S3 <= "00001000";
				S4 <= "00000011";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00000101" => --[1, -6, 125, 11, -4, 1, 0, 0]
				S0 <= "00000001";
				S1 <= "00000110";
				S2 <= "01111101";
				S3 <= "00001011";
				S4 <= "00000100";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00000110" => --[1, -7, 124, 13, -4, 1, 0, 0]
				S0 <= "00000001";
				S1 <= "00000111";
				S2 <= "01111100";
				S3 <= "00001101";
				S4 <= "00000100";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00000111" => --[2, -8, 123, 15, -5, 1, 0, 0]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "01111011";
				S3 <= "00001111";
				S4 <= "00000101";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00001000" => --[2, -9, 122, 18, -6, 1, 0, 0]
				S0 <= "00000010";
				S1 <= "00001001";
				S2 <= "01111010";
				S3 <= "00010010";
				S4 <= "00000110";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00001001" => --[2, -10, 121, 20, -6, 1, 0, 0]
				S0 <= "00000010";
				S1 <= "00001010";
				S2 <= "01111001";
				S3 <= "00010100";
				S4 <= "00000110";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00001010" => --[2, -11, 120, 22, -7, 2, 0, 0]
				S0 <= "00000010";
				S1 <= "00001011";
				S2 <= "01111000";
				S3 <= "00010110";
				S4 <= "00000111";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00001011" => --[2, -12, 119, 25, -8, 2, 0, 0]
				S0 <= "00000010";
				S1 <= "00001100";
				S2 <= "01110111";
				S3 <= "00011001";
				S4 <= "00001000";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00001100" => --[3, -13, 117, 27, -8, 2, 0, 0]
				S0 <= "00000011";
				S1 <= "00001101";
				S2 <= "01110101";
				S3 <= "00011011";
				S4 <= "00001000";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00001101" => --[3, -13, 116, 29, -9, 2, 0, 0]
				S0 <= "00000011";
				S1 <= "00001101";
				S2 <= "01110100";
				S3 <= "00011101";
				S4 <= "00001001";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00001110" => --[3, -14, 114, 32, -10, 3, 0, 0]
				S0 <= "00000011";
				S1 <= "00001110";
				S2 <= "01110010";
				S3 <= "00100000";
				S4 <= "00001010";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00001111" => --[3, -15, 113, 35, -10, 2, 0, 0]
				S0 <= "00000011";
				S1 <= "00001111";
				S2 <= "01110001";
				S3 <= "00100011";
				S4 <= "00001010";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00010000" => --[3, -15, 111, 37, -11, 3, 0, 0]
				S0 <= "00000011";
				S1 <= "00001111";
				S2 <= "01101111";
				S3 <= "00100101";
				S4 <= "00001011";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00010001" => --[3, -16, 109, 40, -11, 3, 0, 0]
				S0 <= "00000011";
				S1 <= "00010000";
				S2 <= "01101101";
				S3 <= "00101000";
				S4 <= "00001011";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00010010" => --[3, -16, 108, 42, -12, 3, 0, 0]
				S0 <= "00000011";
				S1 <= "00010000";
				S2 <= "01101100";
				S3 <= "00101010";
				S4 <= "00001100";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00010011" => --[4, -17, 106, 45, -13, 3, 0, 0]
				S0 <= "00000100";
				S1 <= "00010001";
				S2 <= "01101010";
				S3 <= "00101101";
				S4 <= "00001101";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00010100" => --[4, -17, 104, 47, -13, 3, 0, 0]
				S0 <= "00000100";
				S1 <= "00010001";
				S2 <= "01101000";
				S3 <= "00101111";
				S4 <= "00001101";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00010101" => --[4, -17, 102, 50, -14, 3, 0, 0]
				S0 <= "00000100";
				S1 <= "00010001";
				S2 <= "01100110";
				S3 <= "00110010";
				S4 <= "00001110";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00010110" => --[4, -17, 100, 52, -14, 3, 0, 0]
				S0 <= "00000100";
				S1 <= "00010001";
				S2 <= "01100100";
				S3 <= "00110100";
				S4 <= "00001110";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00010111" => --[4, -18, 98, 55, -15, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01100010";
				S3 <= "00110111";
				S4 <= "00001111";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00011000" => --[4, -18, 96, 58, -15, 3, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01100000";
				S3 <= "00111010";
				S4 <= "00001111";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00011001" => --[4, -18, 94, 60, -16, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01011110";
				S3 <= "00111100";
				S4 <= "00010000";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00011010" => --[4, -18, 91, 63, -16, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01011011";
				S3 <= "00111111";
				S4 <= "00010000";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00011011" => --[4, -18, 89, 65, -16, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01011001";
				S3 <= "01000001";
				S4 <= "00010000";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00011100" => --[4, -18, 87, 68, -17, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01010111";
				S3 <= "01000100";
				S4 <= "00010001";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00011101" => --[4, -18, 85, 70, -17, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01010101";
				S3 <= "01000110";
				S4 <= "00010001";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00011110" => --[4, -18, 82, 73, -17, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01010010";
				S3 <= "01001001";
				S4 <= "00010001";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00011111" => --[4, -18, 80, 75, -17, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01010000";
				S3 <= "01001011";
				S4 <= "00010001";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00100000" => --[4, -18, 78, 78, -18, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010010";
				S2 <= "01001110";
				S3 <= "01001110";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00100001" => --[4, -17, 75, 80, -18, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010001";
				S2 <= "01001011";
				S3 <= "01010000";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00100010" => --[4, -17, 73, 82, -18, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010001";
				S2 <= "01001001";
				S3 <= "01010010";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00100011" => --[4, -17, 70, 85, -18, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010001";
				S2 <= "01000110";
				S3 <= "01010101";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00100100" => --[4, -17, 68, 87, -18, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010001";
				S2 <= "01000100";
				S3 <= "01010111";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00100101" => --[4, -16, 65, 89, -18, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010000";
				S2 <= "01000001";
				S3 <= "01011001";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00100110" => --[4, -16, 63, 91, -18, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010000";
				S2 <= "00111111";
				S3 <= "01011011";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00100111" => --[4, -16, 60, 94, -18, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00010000";
				S2 <= "00111100";
				S3 <= "01011110";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00101000" => --[3, -15, 58, 96, -18, 4, 0, 0]
				S0 <= "00000011";
				S1 <= "00001111";
				S2 <= "00111010";
				S3 <= "01100000";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00101001" => --[4, -15, 55, 98, -18, 4, 0, 0]
				S0 <= "00000100";
				S1 <= "00001111";
				S2 <= "00110111";
				S3 <= "01100010";
				S4 <= "00010010";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00101010" => --[3, -14, 52, 100, -17, 4, 0, 0]
				S0 <= "00000011";
				S1 <= "00001110";
				S2 <= "00110100";
				S3 <= "01100100";
				S4 <= "00010001";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00101011" => --[3, -14, 50, 102, -17, 4, 0, 0]
				S0 <= "00000011";
				S1 <= "00001110";
				S2 <= "00110010";
				S3 <= "01100110";
				S4 <= "00010001";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00101100" => --[3, -13, 47, 104, -17, 4, 0, 0]
				S0 <= "00000011";
				S1 <= "00001101";
				S2 <= "00101111";
				S3 <= "01101000";
				S4 <= "00010001";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00101101" => --[3, -13, 45, 106, -17, 4, 0, 0]
				S0 <= "00000011";
				S1 <= "00001101";
				S2 <= "00101101";
				S3 <= "01101010";
				S4 <= "00010001";
				S5 <= "00000100";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00101110" => --[3, -12, 42, 108, -16, 3, 0, 0]
				S0 <= "00000011";
				S1 <= "00001100";
				S2 <= "00101010";
				S3 <= "01101100";
				S4 <= "00010000";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00101111" => --[3, -11, 40, 109, -16, 3, 0, 0]
				S0 <= "00000011";
				S1 <= "00001011";
				S2 <= "00101000";
				S3 <= "01101101";
				S4 <= "00010000";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00110000" => --[3, -11, 37, 111, -15, 3, 0, 0]
				S0 <= "00000011";
				S1 <= "00001011";
				S2 <= "00100101";
				S3 <= "01101111";
				S4 <= "00001111";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00110001" => --[2, -10, 35, 113, -15, 3, 0, 0]
				S0 <= "00000010";
				S1 <= "00001010";
				S2 <= "00100011";
				S3 <= "01110001";
				S4 <= "00001111";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00110010" => --[3, -10, 32, 114, -14, 3, 0, 0]
				S0 <= "00000011";
				S1 <= "00001010";
				S2 <= "00100000";
				S3 <= "01110010";
				S4 <= "00001110";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00110011" => --[2, -9, 29, 116, -13, 3, 0, 0]
				S0 <= "00000010";
				S1 <= "00001001";
				S2 <= "00011101";
				S3 <= "01110100";
				S4 <= "00001101";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00110100" => --[2, -8, 27, 117, -13, 3, 0, 0]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00011011";
				S3 <= "01110101";
				S4 <= "00001101";
				S5 <= "00000011";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00110101" => --[2, -8, 25, 119, -12, 2, 0, 0]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00011001";
				S3 <= "01110111";
				S4 <= "00001100";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00110110" => --[2, -7, 22, 120, -11, 2, 0, 0]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010110";
				S3 <= "01111000";
				S4 <= "00001011";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00110111" => --[1, -6, 20, 121, -10, 2, 0, 0]
				S0 <= "00000001";
				S1 <= "00000110";
				S2 <= "00010100";
				S3 <= "01111001";
				S4 <= "00001010";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00111000" => --[1, -6, 18, 122, -9, 2, 0, 0]
				S0 <= "00000001";
				S1 <= "00000110";
				S2 <= "00010010";
				S3 <= "01111010";
				S4 <= "00001001";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00111001" => --[1, -5, 15, 123, -8, 2, 0, 0]
				S0 <= "00000001";
				S1 <= "00000101";
				S2 <= "00001111";
				S3 <= "01111011";
				S4 <= "00001000";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00111010" => --[1, -4, 13, 124, -7, 1, 0, 0]
				S0 <= "00000001";
				S1 <= "00000100";
				S2 <= "00001101";
				S3 <= "01111100";
				S4 <= "00000111";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00111011" => --[1, -4, 11, 125, -6, 1, 0, 0]
				S0 <= "00000001";
				S1 <= "00000100";
				S2 <= "00001011";
				S3 <= "01111101";
				S4 <= "00000110";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00111100" => --[1, -3, 8, 126, -5, 1, 0, 0]
				S0 <= "00000001";
				S1 <= "00000011";
				S2 <= "00001000";
				S3 <= "01111110";
				S4 <= "00000101";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00111101" => --[1, -2, 6, 126, -4, 1, 0, 0]
				S0 <= "00000001";
				S1 <= "00000010";
				S2 <= "00000110";
				S3 <= "01111110";
				S4 <= "00000100";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00111110" => --[0, -1, 4, 127, -3, 1, 0, 0]
				S0 <= "00000000";
				S1 <= "00000001";
				S2 <= "00000100";
				S3 <= "01111111";
				S4 <= "00000011";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "00111111" => --[0, 0, 2, 127, -1, 0, 0, 0]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "01111111";
				S4 <= "00000001";
				S5 <= "00000000";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';
				sinalA6 <= '0';

------------------------- Filtro 2------------------------------

			when "01000000" => --[0, 0, 0, 127, 1, 0, 0, 0]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000000";
				S3 <= "01111111";
				S4 <= "00000001";
				S5 <= "00000000";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "01000001" => --[0, 0, -1, 127, 2, 0, 0, 0]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "01111111";
				S4 <= "00000010";
				S5 <= "00000000";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "01000010" => --[0, 1, -3, 127, 4, -2, 1, 0]
				S0 <= "00000000";
				S1 <= "00000001";
				S2 <= "00000011";
				S3 <= "01111111";
				S4 <= "00000100";
				S5 <= "00000010";
				S6 <= "00000001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01000011" => --[0, 1, -5, 127, 6, -2, 1, 0]
				S0 <= "00000000";
				S1 <= "00000001";
				S2 <= "00000101";
				S3 <= "01111111";
				S4 <= "00000110";
				S5 <= "00000010";
				S6 <= "00000001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01000100" => --[0, 2, -6, 126, 8, -3, 1, 0]
				S0 <= "00000000";
				S1 <= "00000010";
				S2 <= "00000110";
				S3 <= "01111110";
				S4 <= "00001000";
				S5 <= "00000011";
				S6 <= "00000001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01000101" => --[-1, 2, -7, 126, 11, -4, 2, -1]
				S0 <= "00000001";
				S1 <= "00000010";
				S2 <= "00000111";
				S3 <= "01111110";
				S4 <= "00001011";
				S5 <= "00000100";
				S6 <= "00000010";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01000110" => --[-1, 3, -8, 125, 13, -5, 2, -1]
				S0 <= "00000001";
				S1 <= "00000011";
				S2 <= "00001000";
				S3 <= "01111101";
				S4 <= "00001101";
				S5 <= "00000101";
				S6 <= "00000010";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01000111" => --[-1, 3, -10, 124, 16, -6, 3, -1]
				S0 <= "00000001";
				S1 <= "00000011";
				S2 <= "00001010";
				S3 <= "01111100";
				S4 <= "00010000";
				S5 <= "00000110";
				S6 <= "00000011";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01001000" => --[-1, 4, -11, 123, 18, -7, 3, -1]
				S0 <= "00000001";
				S1 <= "00000100";
				S2 <= "00001011";
				S3 <= "01111011";
				S4 <= "00010010";
				S5 <= "00000111";
				S6 <= "00000011";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01001001" => --[-1, 4, -12, 122, 20, -7, 3, -1]
				S0 <= "00000001";
				S1 <= "00000100";
				S2 <= "00001100";
				S3 <= "01111010";
				S4 <= "00010100";
				S5 <= "00000111";
				S6 <= "00000011";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01001010" => --[-1, 4, -13, 121, 23, -8, 3, -1]
				S0 <= "00000001";
				S1 <= "00000100";
				S2 <= "00001101";
				S3 <= "01111001";
				S4 <= "00010111";
				S5 <= "00001000";
				S6 <= "00000011";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01001011" => --[-2, 5, -14, 120, 25, -9, 4, -1]
				S0 <= "00000010";
				S1 <= "00000101";
				S2 <= "00001110";
				S3 <= "01111000";
				S4 <= "00011001";
				S5 <= "00001001";
				S6 <= "00000100";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01001100" => --[-1, 5, -15, 119, 27, -10, 4, -1]
				S0 <= "00000001";
				S1 <= "00000101";
				S2 <= "00001111";
				S3 <= "01110111";
				S4 <= "00011011";
				S5 <= "00001010";
				S6 <= "00000100";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01001101" => --[-1, 5, -16, 118, 30, -11, 4, -1]
				S0 <= "00000001";
				S1 <= "00000101";
				S2 <= "00010000";
				S3 <= "01110110";
				S4 <= "00011110";
				S5 <= "00001011";
				S6 <= "00000100";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01001110" => --[-2, 6, -17, 116, 33, -12, 5, -1]
				S0 <= "00000010";
				S1 <= "00000110";
				S2 <= "00010001";
				S3 <= "01110100";
				S4 <= "00100001";
				S5 <= "00001100";
				S6 <= "00000101";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01001111" => --[-2, 6, -17, 114, 35, -12, 5, -1]
				S0 <= "00000010";
				S1 <= "00000110";
				S2 <= "00010001";
				S3 <= "01110010";
				S4 <= "00100011";
				S5 <= "00001100";
				S6 <= "00000101";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01010000" => --[-2, 6, -18, 113, 38, -13, 5, -1]
				S0 <= "00000010";
				S1 <= "00000110";
				S2 <= "00010010";
				S3 <= "01110001";
				S4 <= "00100110";
				S5 <= "00001101";
				S6 <= "00000101";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01010001" => --[-2, 7, -19, 111, 41, -14, 6, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010011";
				S3 <= "01101111";
				S4 <= "00101001";
				S5 <= "00001110";
				S6 <= "00000110";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01010010" => --[-2, 7, -19, 110, 43, -15, 6, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010011";
				S3 <= "01101110";
				S4 <= "00101011";
				S5 <= "00001111";
				S6 <= "00000110";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01010011" => --[-2, 7, -20, 108, 46, -15, 6, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010100";
				S3 <= "01101100";
				S4 <= "00101110";
				S5 <= "00001111";
				S6 <= "00000110";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01010100" => --[-2, 7, -20, 106, 49, -16, 6, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010100";
				S3 <= "01101010";
				S4 <= "00110001";
				S5 <= "00010000";
				S6 <= "00000110";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01010101" => --[-2, 7, -21, 104, 51, -16, 7, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010101";
				S3 <= "01101000";
				S4 <= "00110011";
				S5 <= "00010000";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01010110" => --[-2, 7, -21, 102, 54, -17, 7, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010101";
				S3 <= "01100110";
				S4 <= "00110110";
				S5 <= "00010001";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01010111" => --[-2, 8, -21, 100, 56, -18, 7, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010101";
				S3 <= "01100100";
				S4 <= "00111000";
				S5 <= "00010010";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01011000" => --[-2, 8, -22, 98, 59, -18, 7, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010110";
				S3 <= "01100010";
				S4 <= "00111011";
				S5 <= "00010010";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01011001" => --[-2, 8, -22, 96, 62, -19, 7, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010110";
				S3 <= "01100000";
				S4 <= "00111110";
				S5 <= "00010011";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01011010" => --[-2, 8, -22, 94, 64, -19, 7, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010110";
				S3 <= "01011110";
				S4 <= "01000000";
				S5 <= "00010011";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01011011" => --[-2, 8, -22, 91, 67, -20, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010110";
				S3 <= "01011011";
				S4 <= "01000011";
				S5 <= "00010100";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01011100" => --[-2, 8, -22, 89, 69, -20, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010110";
				S3 <= "01011001";
				S4 <= "01000101";
				S5 <= "00010100";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01011101" => --[-2, 8, -22, 87, 72, -21, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010110";
				S3 <= "01010111";
				S4 <= "01001000";
				S5 <= "00010101";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01011110" => --[-2, 8, -21, 84, 74, -21, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010101";
				S3 <= "01010100";
				S4 <= "01001010";
				S5 <= "00010101";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01011111" => --[-2, 8, -22, 82, 77, -21, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010110";
				S3 <= "01010010";
				S4 <= "01001101";
				S5 <= "00010101";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01100000" => --[-2, 8, -21, 79, 79, -21, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010101";
				S3 <= "01001111";
				S4 <= "01001111";
				S5 <= "00010101";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01100001" => --[-2, 8, -21, 77, 82, -22, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010101";
				S3 <= "01001101";
				S4 <= "01010010";
				S5 <= "00010110";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01100010" => --[-2, 8, -21, 74, 84, -21, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010101";
				S3 <= "01001010";
				S4 <= "01010100";
				S5 <= "00010101";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01100011" => --[-2, 8, -21, 72, 87, -22, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010101";
				S3 <= "01001000";
				S4 <= "01010111";
				S5 <= "00010110";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01100100" => --[-2, 8, -20, 69, 89, -22, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010100";
				S3 <= "01000101";
				S4 <= "01011001";
				S5 <= "00010110";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01100101" => --[-2, 8, -20, 67, 91, -22, 8, -2]
				S0 <= "00000010";
				S1 <= "00001000";
				S2 <= "00010100";
				S3 <= "01000011";
				S4 <= "01011011";
				S5 <= "00010110";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01100110" => --[-2, 7, -19, 64, 94, -22, 8, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010011";
				S3 <= "01000000";
				S4 <= "01011110";
				S5 <= "00010110";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01100111" => --[-2, 7, -19, 62, 96, -22, 8, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010011";
				S3 <= "00111110";
				S4 <= "01100000";
				S5 <= "00010110";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01101000" => --[-2, 7, -18, 59, 98, -22, 8, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010010";
				S3 <= "00111011";
				S4 <= "01100010";
				S5 <= "00010110";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01101001" => --[-2, 7, -18, 56, 100, -21, 8, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010010";
				S3 <= "00111000";
				S4 <= "01100100";
				S5 <= "00010101";
				S6 <= "00001000";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01101010" => --[-2, 7, -17, 54, 102, -21, 7, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010001";
				S3 <= "00110110";
				S4 <= "01100110";
				S5 <= "00010101";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01101011" => --[-2, 7, -16, 51, 104, -21, 7, -2]
				S0 <= "00000010";
				S1 <= "00000111";
				S2 <= "00010000";
				S3 <= "00110011";
				S4 <= "01101000";
				S5 <= "00010101";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01101100" => --[-2, 6, -16, 49, 106, -20, 7, -2]
				S0 <= "00000010";
				S1 <= "00000110";
				S2 <= "00010000";
				S3 <= "00110001";
				S4 <= "01101010";
				S5 <= "00010100";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01101101" => --[-2, 6, -15, 46, 108, -20, 7, -2]
				S0 <= "00000010";
				S1 <= "00000110";
				S2 <= "00001111";
				S3 <= "00101110";
				S4 <= "01101100";
				S5 <= "00010100";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01101110" => --[-2, 6, -15, 43, 110, -19, 7, -2]
				S0 <= "00000010";
				S1 <= "00000110";
				S2 <= "00001111";
				S3 <= "00101011";
				S4 <= "01101110";
				S5 <= "00010011";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01101111" => --[-2, 6, -14, 41, 111, -19, 7, -2]
				S0 <= "00000010";
				S1 <= "00000110";
				S2 <= "00001110";
				S3 <= "00101001";
				S4 <= "01101111";
				S5 <= "00010011";
				S6 <= "00000111";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01110000" => --[-1, 5, -13, 38, 113, -18, 6, -2]
				S0 <= "00000001";
				S1 <= "00000101";
				S2 <= "00001101";
				S3 <= "00100110";
				S4 <= "01110001";
				S5 <= "00010010";
				S6 <= "00000110";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01110001" => --[-1, 5, -12, 35, 114, -17, 6, -2]
				S0 <= "00000001";
				S1 <= "00000101";
				S2 <= "00001100";
				S3 <= "00100011";
				S4 <= "01110010";
				S5 <= "00010001";
				S6 <= "00000110";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01110010" => --[-1, 5, -12, 33, 116, -17, 6, -2]
				S0 <= "00000001";
				S1 <= "00000101";
				S2 <= "00001100";
				S3 <= "00100001";
				S4 <= "01110100";
				S5 <= "00010001";
				S6 <= "00000110";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01110011" => --[-1, 4, -11, 30, 118, -16, 5, -1]
				S0 <= "00000001";
				S1 <= "00000100";
				S2 <= "00001011";
				S3 <= "00011110";
				S4 <= "01110110";
				S5 <= "00010000";
				S6 <= "00000101";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01110100" => --[-1, 4, -10, 27, 119, -15, 5, -1]
				S0 <= "00000001";
				S1 <= "00000100";
				S2 <= "00001010";
				S3 <= "00011011";
				S4 <= "01110111";
				S5 <= "00001111";
				S6 <= "00000101";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01110101" => --[-1, 4, -9, 25, 120, -14, 5, -2]
				S0 <= "00000001";
				S1 <= "00000100";
				S2 <= "00001001";
				S3 <= "00011001";
				S4 <= "01111000";
				S5 <= "00001110";
				S6 <= "00000101";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01110110" => --[-1, 3, -8, 23, 121, -13, 4, -1]
				S0 <= "00000001";
				S1 <= "00000011";
				S2 <= "00001000";
				S3 <= "00010111";
				S4 <= "01111001";
				S5 <= "00001101";
				S6 <= "00000100";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01110111" => --[-1, 3, -7, 20, 122, -12, 4, -1]
				S0 <= "00000001";
				S1 <= "00000011";
				S2 <= "00000111";
				S3 <= "00010100";
				S4 <= "01111010";
				S5 <= "00001100";
				S6 <= "00000100";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01111000" => --[-1, 3, -7, 18, 123, -11, 4, -1]
				S0 <= "00000001";
				S1 <= "00000011";
				S2 <= "00000111";
				S3 <= "00010010";
				S4 <= "01111011";
				S5 <= "00001011";
				S6 <= "00000100";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01111001" => --[-1, 3, -6, 16, 124, -10, 3, -1]
				S0 <= "00000001";
				S1 <= "00000011";
				S2 <= "00000110";
				S3 <= "00010000";
				S4 <= "01111100";
				S5 <= "00001010";
				S6 <= "00000011";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01111010" => --[-1, 2, -5, 13, 125, -8, 3, -1]
				S0 <= "00000001";
				S1 <= "00000010";
				S2 <= "00000101";
				S3 <= "00001101";
				S4 <= "01111101";
				S5 <= "00001000";
				S6 <= "00000011";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01111011" => --[-1, 2, -4, 11, 126, -7, 2, -1]
				S0 <= "00000001";
				S1 <= "00000010";
				S2 <= "00000100";
				S3 <= "00001011";
				S4 <= "01111110";
				S5 <= "00000111";
				S6 <= "00000010";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01111100" => --[0, 1, -3, 8, 126, -6, 2, 0]
				S0 <= "00000000";
				S1 <= "00000001";
				S2 <= "00000011";
				S3 <= "00001000";
				S4 <= "01111110";
				S5 <= "00000110";
				S6 <= "00000010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01111101" => --[0, 1, -2, 6, 127, -5, 1, 0]
				S0 <= "00000000";
				S1 <= "00000001";
				S2 <= "00000010";
				S3 <= "00000110";
				S4 <= "01111111";
				S5 <= "00000101";
				S6 <= "00000001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01111110" => --[0, 1, -2, 4, 127, -3, 1, 0]
				S0 <= "00000000";
				S1 <= "00000001";
				S2 <= "00000010";
				S3 <= "00000100";
				S4 <= "01111111";
				S5 <= "00000011";
				S6 <= "00000001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '1';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

			when "01111111" => --[0, 0, 0, 2, 127, -1, 0, 0]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000000";
				S3 <= "00000010";
				S4 <= "01111111";
				S5 <= "00000001";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
				sinalA6 <= '0';

------------------------- Filtro 3------------------------------

			when "10000000" => --[0, 0, 0, 1, 127, 0, 0, 0]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000000";
				S3 <= "00000001";
				S4 <= "01111111";
				S5 <= "00000000";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "10000001" => --[0, 0, 0, -1, 127, 2, 0, 0]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000000";
				S3 <= "00000001";
				S4 <= "01111111";
				S5 <= "00000010";
				S6 <= "00000000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '0';

			when "10000010" => --[0, 0, 1, -3, 127, 4, -1, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000011";
				S4 <= "01111111";
				S5 <= "00000100";
				S6 <= "00000001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10000011" => --[0, 0, 1, -4, 126, 6, -2, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000100";
				S4 <= "01111110";
				S5 <= "00000110";
				S6 <= "00000010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10000100" => --[0, 0, 1, -5, 126, 8, -3, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000101";
				S4 <= "01111110";
				S5 <= "00001000";
				S6 <= "00000011";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10000101" => --[0, 0, 1, -6, 125, 11, -4, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000110";
				S4 <= "01111101";
				S5 <= "00001011";
				S6 <= "00000100";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10000110" => --[0, 0, 1, -7, 124, 13, -4, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000111";
				S4 <= "01111100";
				S5 <= "00001101";
				S6 <= "00000100";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10000111" => --[0, 0, 2, -8, 123, 15, -5, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00001000";
				S4 <= "01111011";
				S5 <= "00001111";
				S6 <= "00000101";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10001000" => --[0, 0, 2, -9, 122, 18, -6, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00001001";
				S4 <= "01111010";
				S5 <= "00010010";
				S6 <= "00000110";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10001001" => --[0, 0, 2, -10, 121, 20, -6, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00001010";
				S4 <= "01111001";
				S5 <= "00010100";
				S6 <= "00000110";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10001010" => --[0, 0, 2, -11, 120, 22, -7, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00001011";
				S4 <= "01111000";
				S5 <= "00010110";
				S6 <= "00000111";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10001011" => --[0, 0, 2, -12, 119, 25, -8, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00001100";
				S4 <= "01110111";
				S5 <= "00011001";
				S6 <= "00001000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10001100" => --[0, 0, 3, -13, 117, 27, -8, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001101";
				S4 <= "01110101";
				S5 <= "00011011";
				S6 <= "00001000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10001101" => --[0, 0, 3, -13, 116, 29, -9, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001101";
				S4 <= "01110100";
				S5 <= "00011101";
				S6 <= "00001001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10001110" => --[0, 0, 3, -14, 114, 32, -10, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001110";
				S4 <= "01110010";
				S5 <= "00100000";
				S6 <= "00001010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10001111" => --[0, 0, 3, -15, 113, 35, -10, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001111";
				S4 <= "01110001";
				S5 <= "00100011";
				S6 <= "00001010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10010000" => --[0, 0, 3, -15, 111, 37, -11, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001111";
				S4 <= "01101111";
				S5 <= "00100101";
				S6 <= "00001011";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10010001" => --[0, 0, 3, -16, 109, 40, -11, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00010000";
				S4 <= "01101101";
				S5 <= "00101000";
				S6 <= "00001011";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10010010" => --[0, 0, 3, -16, 108, 42, -12, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00010000";
				S4 <= "01101100";
				S5 <= "00101010";
				S6 <= "00001100";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10010011" => --[0, 0, 4, -17, 106, 45, -13, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010001";
				S4 <= "01101010";
				S5 <= "00101101";
				S6 <= "00001101";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10010100" => --[0, 0, 4, -17, 104, 47, -13, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010001";
				S4 <= "01101000";
				S5 <= "00101111";
				S6 <= "00001101";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10010101" => --[0, 0, 4, -17, 102, 50, -14, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010001";
				S4 <= "01100110";
				S5 <= "00110010";
				S6 <= "00001110";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10010110" => --[0, 0, 4, -17, 100, 52, -14, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010001";
				S4 <= "01100100";
				S5 <= "00110100";
				S6 <= "00001110";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10010111" => --[0, 0, 4, -18, 98, 55, -15, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01100010";
				S5 <= "00110111";
				S6 <= "00001111";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10011000" => --[0, 0, 4, -18, 96, 58, -15, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01100000";
				S5 <= "00111010";
				S6 <= "00001111";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10011001" => --[0, 0, 4, -18, 94, 60, -16, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01011110";
				S5 <= "00111100";
				S6 <= "00010000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10011010" => --[0, 0, 4, -18, 91, 63, -16, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01011011";
				S5 <= "00111111";
				S6 <= "00010000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10011011" => --[0, 0, 4, -18, 89, 65, -16, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01011001";
				S5 <= "01000001";
				S6 <= "00010000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10011100" => --[0, 0, 4, -18, 87, 68, -17, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01010111";
				S5 <= "01000100";
				S6 <= "00010001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10011101" => --[0, 0, 4, -18, 85, 70, -17, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01010101";
				S5 <= "01000110";
				S6 <= "00010001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10011110" => --[0, 0, 4, -18, 82, 73, -17, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01010010";
				S5 <= "01001001";
				S6 <= "00010001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10011111" => --[0, 0, 4, -18, 80, 75, -17, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01010000";
				S5 <= "01001011";
				S6 <= "00010001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10100000" => --[0, 0, 4, -18, 78, 78, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010010";
				S4 <= "01001110";
				S5 <= "01001110";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10100001" => --[0, 0, 4, -17, 75, 80, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010001";
				S4 <= "01001011";
				S5 <= "01010000";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10100010" => --[0, 0, 4, -17, 73, 82, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010001";
				S4 <= "01001001";
				S5 <= "01010010";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10100011" => --[0, 0, 4, -17, 70, 85, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010001";
				S4 <= "01000110";
				S5 <= "01010101";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10100100" => --[0, 0, 4, -17, 68, 87, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010001";
				S4 <= "01000100";
				S5 <= "01010111";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10100101" => --[0, 0, 4, -16, 65, 89, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010000";
				S4 <= "01000001";
				S5 <= "01011001";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10100110" => --[0, 0, 4, -16, 63, 91, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010000";
				S4 <= "00111111";
				S5 <= "01011011";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10100111" => --[0, 0, 4, -16, 60, 84, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00010000";
				S4 <= "00111100";
				S5 <= "01010100";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10101000" => --[0, 0, 3, -15, 58, 96, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001111";
				S4 <= "00111010";
				S5 <= "01100000";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10101001" => --[0, 0, 4, -15, 55, 98, -18, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000100";
				S3 <= "00001111";
				S4 <= "00110111";
				S5 <= "01100010";
				S6 <= "00010010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10101010" => --[0, 0, 3, -14, 52, 100, -17, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001110";
				S4 <= "00110100";
				S5 <= "01100100";
				S6 <= "00010001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10101011" => --[0, 0, 3, -14, 50, 102, -17, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001110";
				S4 <= "00110010";
				S5 <= "01100110";
				S6 <= "00010001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10101100" => --[0, 0, 3, -13, 47, 104, -17, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001101";
				S4 <= "00101111";
				S5 <= "01101000";
				S6 <= "00010001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10101101" => --[0, 0, 3, -13, 45, 106, -17, 4]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001101";
				S4 <= "00101101";
				S5 <= "01101010";
				S6 <= "00010001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10101110" => --[0, 0, 3, -12, 42, 108, -16, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001100";
				S4 <= "00101010";
				S5 <= "01101100";
				S6 <= "00010000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10101111" => --[0, 0, 3, -11, 40, 109, -16, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001011";
				S4 <= "00101000";
				S5 <= "01101101";
				S6 <= "00010000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10110000" => --[0, 0, 3, -11, 37, 111, -15, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001011";
				S4 <= "00100101";
				S5 <= "01101111";
				S6 <= "00001111";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10110001" => --[0, 0, 2, -10, 35, 113, -15, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00001010";
				S4 <= "00100011";
				S5 <= "01110001";
				S6 <= "00001111";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10110010" => --[0, 0, 3, -10, 32, 114, -14, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000011";
				S3 <= "00001010";
				S4 <= "00100000";
				S5 <= "01110010";
				S6 <= "00001110";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10110011" => --[0, 0, 2, -9, 29, 116, -13, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00001001";
				S4 <= "00011101";
				S5 <= "01110100";
				S6 <= "00001101";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10110100" => --[0, 0, 2, -8, 27, 117, -13, 3]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00001000";
				S4 <= "00011011";
				S5 <= "01110101";
				S6 <= "00001101";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10110101" => --[0, 0, 2, -8, 25, 119, -12, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00001000";
				S4 <= "00011001";
				S5 <= "01110111";
				S6 <= "00001100";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10110110" => --[0, 0, 2, -7, 22, 120, -11, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000010";
				S3 <= "00000111";
				S4 <= "00010110";
				S5 <= "01111000";
				S6 <= "00001011";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10110111" => --[0, 0, 1, -6, 20, 121, -10, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000110";
				S4 <= "00010100";
				S5 <= "01111001";
				S6 <= "00001010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10111000" => --[0, 0, 1, -6, 18, 122, -9, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000110";
				S4 <= "00010010";
				S5 <= "01111010";
				S6 <= "00001001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10111001" => --[0, 0, 1, -5, 15, 123, -8, 2]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000101";
				S4 <= "00001111";
				S5 <= "01111011";
				S6 <= "00001000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10111010" => --[0, 0, 1, -4, 13, 124, -7, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000100";
				S4 <= "00001101";
				S5 <= "01111100";
				S6 <= "00000111";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10111011" => --[0, 0, 1, -4, 11, 125, -6, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000100";
				S4 <= "00001011";
				S5 <= "01111101";
				S6 <= "00000110";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10111100" => --[0, 0, 1, -3, 8, 126, -5, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000011";
				S4 <= "00001000";
				S5 <= "01111110";
				S6 <= "00000101";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10111101" => --[0, 0, 1, -2, 6, 126, -4, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000001";
				S3 <= "00000010";
				S4 <= "00000110";
				S5 <= "01111110";
				S6 <= "00000100";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10111110" => --[0, 0, 0, -1, 4, 127, -3, 1]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000000";
				S3 <= "00000001";
				S4 <= "00000100";
				S5 <= "01111111";
				S6 <= "00000011";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when "10111111" => --[0, 0, 0, 0, 2, 127, -1, 0]
				S0 <= "00000000";
				S1 <= "00000000";
				S2 <= "00000000";
				S3 <= "00000000";
				S4 <= "00000010";
				S5 <= "01111111";
				S6 <= "00000001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA2 <= '0';
				sinalA3 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
				sinalA6 <= '1';

			when others =>
				aux8 <= "00";
		
		end case;

	end process;

end comportamento;