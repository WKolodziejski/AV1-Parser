library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_signed.all;
use ieee.numeric_std.all; 

entity Escolha is
	port(vet_sel: in std_logic_vector(7 downto 0);
		S0, S3: out std_logic_vector(2 downto 0);
		S1, S2: out std_logic_vector(5 downto 0);
		sinalA0, sinalA1: out std_logic
		);
end Escolha;


architecture comportamento of Escolha is
	signal aux8: signed (1 downto 0);
	begin
	process (vet_sel)
	begin

		case vet_sel is


------------------------- Filtro 1------------------------------

			when "00000000" => --[0, 0, 128, 0, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "001001";
				S3 <= "001001";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00000001" => --[2, -4, 108, 16, 4, 2]
				S0 <= "001";
				S1 <= "010";
				S2 <= "000111";
				S3 <= "000001";
				S4 <= "010";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00000010" => --[4, -16, 108, 44, -16, 4]
				S0 <= "010";
				S1 <= "100";
				S2 <= "000111";
				S3 <= "000100";
				S4 <= "100";
				S5 <= "010";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00000011" => --[2, -16, 84, 64, -8, 2]
				S0 <= "001";
				S1 <= "100";
				S2 <= "000110";
				S3 <= "000101";
				S4 <= "011";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00000100" => --[4, -32, 84, 84, -16, 4]
				S0 <= "010";
				S1 <= "101";
				S2 <= "000110";
				S3 <= "000110";
				S4 <= "100";
				S5 <= "010";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00000101" => --[2, -8, 64, 84, -16, 2]
				S0 <= "001";
				S1 <= "011";
				S2 <= "000101";
				S3 <= "000110";
				S4 <= "100";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00000110" => --[4, -16, 44, 108, -16, 4]
				S0 <= "010";
				S1 <= "100";
				S2 <= "000100";
				S3 <= "000111";
				S4 <= "100";
				S5 <= "010";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00000111" => --[2, 4, 16, 108, -4, 2]
				S0 <= "001";
				S1 <= "010";
				S2 <= "000001";
				S3 <= "000111";
				S4 <= "010";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '1';
				sinalA5 <= '0';

------------------------- Filtro 2------------------------------

			when "00001000" => --[0, 0, 128, 0, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "001001";
				S3 <= "001001";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00001001" => --[2, 32, 64, 20, 8, 2]
				S0 <= "001";
				S1 <= "101";
				S2 <= "000101";
				S3 <= "000010";
				S4 <= "011";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00001010" => --[-2, 32, 64, 32, 4, -2]
				S0 <= "001";
				S1 <= "101";
				S2 <= "000101";
				S3 <= "000011";
				S4 <= "010";
				S5 <= "001";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
			when "00001011" => --[2, 32, 44, 32, 16, 2]
				S0 <= "001";
				S1 <= "101";
				S2 <= "000100";
				S3 <= "000011";
				S4 <= "100";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00001100" => --[4, 16, 44, 44, 16, 4]
				S0 <= "010";
				S1 <= "100";
				S2 <= "000100";
				S3 <= "000100";
				S4 <= "100";
				S5 <= "010";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00001101" => --[2, 16, 32, 44, 32, 2]
				S0 <= "001";
				S1 <= "100";
				S2 <= "000011";
				S3 <= "000100";
				S4 <= "101";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00001110" => --[-2, 4, 32, 64, 32, -2]
				S0 <= "001";
				S1 <= "010";
				S2 <= "000011";
				S3 <= "000101";
				S4 <= "101";
				S5 <= "001";
				sinalA0 <= '1';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '1';
			when "00001111" => --[2, 8, 20, 64, 32, 2]
				S0 <= "001";
				S1 <= "011";
				S2 <= "000010";
				S3 <= "000101";
				S4 <= "101";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';

------------------------- Filtro 3------------------------------

			when "00010000" => --[0, 0, 128, 0, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "001001";
				S3 <= "001001";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00010001" => --[4, -2, 108, 16, -2, 4]
				S0 <= "010";
				S1 <= "001";
				S2 <= "000111";
				S3 <= "000001";
				S4 <= "001";
				S5 <= "010";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00010010" => --[4, -16, 108, 44, -16, 4]
				S0 <= "010";
				S1 <= "100";
				S2 <= "000111";
				S3 <= "000100";
				S4 <= "100";
				S5 <= "010";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00010011" => --[2, -32, 108, 64, -16, 2]
				S0 <= "001";
				S1 <= "101";
				S2 <= "000111";
				S3 <= "000101";
				S4 <= "100";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00010100" => --[4, -32, 84, 84, -16, 4]
				S0 <= "010";
				S1 <= "101";
				S2 <= "000110";
				S3 <= "000110";
				S4 <= "100";
				S5 <= "010";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00010101" => --[2, -16, 64, 108, -32, 2]
				S0 <= "001";
				S1 <= "100";
				S2 <= "000101";
				S3 <= "000111";
				S4 <= "101";
				S5 <= "001";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00010110" => --[4, -16, 44, 108, -16, 4]
				S0 <= "010";
				S1 <= "100";
				S2 <= "000100";
				S3 <= "000111";
				S4 <= "100";
				S5 <= "010";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00010111" => --[4, -2, 16, 108, -2, 4]
				S0 <= "010";
				S1 <= "001";
				S2 <= "000001";
				S3 <= "000111";
				S4 <= "001";
				S5 <= "010";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';

------------------------- Filtro 4------------------------------

			when "00011000" => --[0, 0, 128, 0, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "001001";
				S3 <= "001001";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00011001" => --[0, 0, 108, 20, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "000111";
				S3 <= "000010";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00011010" => --[0, 0, 108, 20, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "000111";
				S3 <= "000010";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00011011" => --[0, 0, 84, 44, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "000110";
				S3 <= "000100";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00011100" => --[0, 0, 64, 64, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "000101";
				S3 <= "000101";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00011101" => --[0, 0, 44, 84, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "000100";
				S3 <= "000110";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00011110" => --[0, 0, 20, 108, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "000010";
				S3 <= "000111";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00011111" => --[0, 0, 20, 108, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "000010";
				S3 <= "000111";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';

------------------------- Filtro 5------------------------------

			when "00100000" => --[0, 0, 128, 0, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "001001";
				S3 <= "001001";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00100001" => --[0, 2, 108, 16, 2, 0]
				S0 <= "000";
				S1 <= "001";
				S2 <= "000111";
				S3 <= "000001";
				S4 <= "001";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00100010" => --[0, -16, 108, 44, -8, 0]
				S0 <= "000";
				S1 <= "100";
				S2 <= "000111";
				S3 <= "000100";
				S4 <= "011";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00100011" => --[0, -16, 84, 64, -4, 0]
				S0 <= "000";
				S1 <= "100";
				S2 <= "000110";
				S3 <= "000101";
				S4 <= "010";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00100100" => --[0, -32, 84, 84, -8, 0]
				S0 <= "000";
				S1 <= "101";
				S2 <= "000110";
				S3 <= "000110";
				S4 <= "011";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00100101" => --[0, -4, 64, 84, -16, 0]
				S0 <= "000";
				S1 <= "010";
				S2 <= "000101";
				S3 <= "000110";
				S4 <= "100";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00100110" => --[0, -8, 44, 108, -16, 0]
				S0 <= "000";
				S1 <= "011";
				S2 <= "000100";
				S3 <= "000111";
				S4 <= "100";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '1';
				sinalA4 <= '1';
				sinalA5 <= '0';
			when "00100111" => --[0, 2, 16, 108, 2, 0]
				S0 <= "000";
				S1 <= "001";
				S2 <= "000001";
				S3 <= "000111";
				S4 <= "001";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';

------------------------- Filtro 6------------------------------

			when "00101000" => --[0, 0, 128, 0, 0, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "001001";
				S3 <= "001001";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00101001" => --[0, 32, 64, 32, 0, 0]
				S0 <= "000";
				S1 <= "101";
				S2 <= "000101";
				S3 <= "000011";
				S4 <= "000";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00101010" => --[0, 16, 64, 44, 4, 0]
				S0 <= "000";
				S1 <= "100";
				S2 <= "000101";
				S3 <= "000100";
				S4 <= "010";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00101011" => --[0, 16, 64, 44, 4, 0]
				S0 <= "000";
				S1 <= "100";
				S2 <= "000101";
				S3 <= "000100";
				S4 <= "010";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00101100" => --[0, 32, 44, 44, 8, 0]
				S0 <= "000";
				S1 <= "101";
				S2 <= "000100";
				S3 <= "000100";
				S4 <= "011";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00101101" => --[0, 4, 44, 64, 16, 0]
				S0 <= "000";
				S1 <= "010";
				S2 <= "000100";
				S3 <= "000101";
				S4 <= "100";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00101110" => --[0, 4, 44, 64, 16, 0]
				S0 <= "000";
				S1 <= "010";
				S2 <= "000100";
				S3 <= "000101";
				S4 <= "100";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when "00101111" => --[0, 0, 32, 64, 32, 0]
				S0 <= "000";
				S1 <= "000";
				S2 <= "000011";
				S3 <= "000101";
				S4 <= "101";
				S5 <= "000";
				sinalA0 <= '0';
				sinalA1 <= '0';
				sinalA4 <= '0';
				sinalA5 <= '0';
			when others =>
				aux8 <= "00";
		
		end case;

	end process;

end comportamento;